-- Cardbus MIMO1 Wireless Com Features
  constant CFG_CMIMO1_ENABLE : integer := CONFIG_CMIMO1_ENABLE;
  constant CFG_CMIMO1_IO : integer := 16#CONFIG_CMIMO1_IO#;
  constant CFG_CMIMO1_RFCTRL_IO_OFFSET : integer := 16#CONFIG_CMIMO1_RFCTRL_IO_OFFSET#;
  constant CFG_CMIMO1_ADAC_IO_OFFSET : integer := 16#CONFIG_CMIMO1_ADAC_IO_OFFSET#;
  constant CFG_CMIMO1_SPI_IO_OFFSET : integer := 16#CONFIG_CMIMO1_SPI_IO_OFFSET#;
  constant CFG_CMIMO1_IDROMEL_SPI_IO_OFFSET : integer := 16#CONFIG_CMIMO1_IDROMEL_SPI_IO_OFFSET#;
  constant CFG_CMIMO1_HADDR : integer := 16#CONFIG_CMIMO1_HADDR#;
  constant CFG_CMIMO1_HMASK : integer := 16#CONFIG_CMIMO1_HMASK#;
  constant CFG_CMIMO1_ADAC_ADC0_HOFFSET : integer := 16#CONFIG_CMIMO1_ADAC_ADC0_HOFFSET#;
  constant CFG_CMIMO1_ADAC_RAMADC0_KBSZ : integer := CONFIG_CMIMO1_ADAC_RAMADC0_KBSZ;
  constant CFG_CMIMO1_ADAC_ADC1_HOFFSET : integer := 16#CONFIG_CMIMO1_ADAC_ADC1_HOFFSET#;
  constant CFG_CMIMO1_ADAC_RAMADC1_KBSZ : integer := CONFIG_CMIMO1_ADAC_RAMADC1_KBSZ;
  constant CFG_CMIMO1_ADAC_DAC0_HOFFSET : integer := 16#CONFIG_CMIMO1_ADAC_DAC0_HOFFSET#;
  constant CFG_CMIMO1_ADAC_RAMDAC0_KBSZ : integer := CONFIG_CMIMO1_ADAC_RAMDAC0_KBSZ;
  constant CFG_CMIMO1_ADAC_DAC1_HOFFSET : integer := 16#CONFIG_CMIMO1_ADAC_DAC1_HOFFSET#;
  constant CFG_CMIMO1_ADAC_RAMDAC1_KBSZ : integer := CONFIG_CMIMO1_ADAC_RAMDAC1_KBSZ;
  constant CFG_CMIMO1_IRQ : integer := CONFIG_CMIMO1_IRQ;

